`timescale 1ns / 1ps

module bcd_2dec(
    input clk,
    input rst,
    input up,
    input cnten1,
    input cnten2,
    output [3:0] bcd0,
    output [3:0] bcd1
    );


endmodule
